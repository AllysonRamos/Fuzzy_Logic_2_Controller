module compara_Maximo  (A,B,S);

input [7:0] A,B;

output [7:0] S;

assign S =(A>B)?A:B;

endmodule
